module exec
#(
    parameter M_WIDTH = 8,
    parameter OP_LUI = 7'b0110111,
    parameter OP_AIUPC = 7'b0010111,
    parameter OP_JAL = 7'b1101111,
    parameter OP_JALR = 7'b1100111,
    parameter OP_LOAD = 7'b0000011,
    parameter OP_STORE = 7'b0100011,
    parameter OP_BRANCH = 7'b1100011,
    parameter OP_INTEGER_IMM = 7'b0010011,
    parameter OP_INTEGER = 7'b0110011
)
(
    input en,
    input clk,
    input [3:0] op,
    input [6:0] funct7,
    input [2:0] funct3,
    input [M_WIDTH-1:0] pc_in,
    input [M_WIDTH-1:0] rs1,
    input [M_WIDTH-1:0] rs2,
    input [M_WIDTH-1:0] imm,
    input [M_WIDTH-1:0] mem_data_in,
    input mem_ready,
    output reg [M_WIDTH-1:0] pc_out,
    output reg [M_WIDTH-1:0] val_out,
    output reg [M_WIDTH-1:0] mem_addr,
    output reg [M_WIDTH-1:0] mem_data_out,
    output reg mem_req,
    output reg mem_we,
    output reg flush_pipeline,
    output reg ready
);

reg [1:0] cycle;

wire [M_WIDTH-1:0] imm_pl_rs1, next_pc;

assign imm_pl_rs1 = imm + rs1;
assign next_pc = pc_in + 4;

always @ (posedge clk) begin
    if (en) begin
        if (op == OP_LOAD || op == OP_STORE) begin
            ready <= cycle == 2;

            if (cycle == 0) begin
                mem_addr <= imm_pl_rs1;
                mem_we <= op == OP_STORE;
                mem_data_out <= rs2;
                mem_req <= 1;
                cycle <= 1;
            end

            if (cycle == 1 && mem_ready) begin
                cycle <= 2;
                mem_req <= 0;
                val_out <= mem_data_in;
            end
        end

        else begin
            ready <= cycle;
            if (cycle == 0) begin
                casez (op)
                    OP_LUI: val_out <= imm;
                    OP_AIUPC: val_out <= pc_in + imm;
                    OP_JAL: begin
                        pc_out <= pc_in + imm;
                        val_out <= next_pc;
                        flush_pipeline <= 1;
                    end
                    OP_JALR: begin
                        pc_out <= {imm_pl_rs1[M_WIDTH-1:1], 1'b0};
                        val_out <= next_pc;
                        flush_pipeline <= 1;
                    end
                    OP_INTEGER_IMM: begin
                        case (funct3)
                            0: val_out <= imm_pl_rs1;
                            1: val_out <= rs1 << imm[4:0];
                            2: val_out <= rs1 < imm;
                            3: val_out <= {1'b0, rs1} < {1'b0, imm};
                            4: val_out <= rs1 ^ imm;
                            5: val_out <= imm[30] ? rs1 >>> imm[4:0] : rs1 >> imm[4:0];
                            6: val_out <= rs1 | imm;
                            7: val_out <= rs1 & imm;
                        endcase
                    end
                    OP_INTEGER: begin
                        case (funct3)
                            0: val_out <= rs1 + rs2;
                            1: val_out <= rs1 << rs2;
                            2: val_out <= rs1 < rs2;
                            3: val_out <= {1'b0, rs1} < {1'b0, rs2};
                            4: val_out <= rs1 ^ rs2;
                            5: val_out <= funct7[5] ? rs1 >>> rs2 : rs1 >> rs2;
                            6: val_out <= rs1 | rs2;
                            7: val_out <= rs1 & rs2;
                        endcase
                    end
                endcase
                cycle <= 1;
            end
        end
    end else begin
        ready <= 0;
        cycle <= 0;
        mem_req <= 0;
        flush_pipeline <= 0;
    end
end

endmodule
